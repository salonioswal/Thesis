library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all;
use work.my_package.all; 
use work.all;


ENTITY ROM_weights is 
PORT ( rd_addr : in unsigned (7 downto 0);
       data_out: out signed (data_width-1 downto 0));
END ROM_weights;

ARCHITECTURE behavior OF ROM_weights IS 
signal all_coeffs: RF(255 downto 0);
begin
      all_coeffs(0) <= signed(13,data_width);
      all_coeffs(1) <= signed(15,data_width);
      all_coeffs(2) <= signed(13,data_width);
      all_coeffs(3) <= signed(0,data_width);
      all_coeffs(4) <= signed(2,data_width);
      all_coeffs(5) <= signed(7,data_width);
      all_coeffs(6) <= signed(8,data_width);
      all_coeffs(7) <= signed(4,data_width);
      all_coeffs(8) <= signed(6,data_width);
      all_coeffs(9) <= signed(5,data_width);
      all_coeffs(10)<=signed(3,data_width);
      all_coeffs(11) <= signed(14,data_width);
      all_coeffs(12) <= signed(15,data_width);
      all_coeffs(13) <= signed(14,data_width);
      all_coeffs(14) <= signed(1,data_width);
      all_coeffs(15) <= signed(7,data_width);
      all_coeffs(16) <= signed(15,data_width);
      all_coeffs(17) <= signed(2,data_width);
      all_coeffs(18) <= signed(9,data_width);
      all_coeffs(19) <= signed(9,data_width);
      all_coeffs(20) <= signed(2,data_width);
      all_coeffs(21)<= signed(2,data_width);
      all_coeffs(22) <= signed(2,data_width);
      all_coeffs(23) <= signed(7,data_width);
      all_coeffs(24) <= signed(10,data_width);
      all_coeffs(25) <= signed(13,data_width);
      all_coeffs(26) <= signed(7,data_width);
      all_coeffs(27) <= signed(5,data_width);
      all_coeffs(28) <= signed(2,data_width);
      all_coeffs(29) <= signed(7,data_width);
      all_coeffs(30) <= signed(1,data_width);
      all_coeffs(31) <= signed(12,data_width);
      all_coeffs(32) <= signed(6,data_width);
      all_coeffs(33) <= signed(14,data_width);
      all_coeffs(34) <= signed(12,data_width);
      all_coeffs(35) <= signed(12,data_width);
      all_coeffs(36) <= signed(11,data_width);
      all_coeffs(37) <= signed(10,data_width);
      all_coeffs(38) <= signed(9,data_width);
      all_coeffs(39) <= signed(4,data_width);
      all_coeffs(40) <= signed(5,data_width);
      all_coeffs(41) <= signed(0,data_width);
      all_coeffs(42) <= signed(4,data_width);
      all_coeffs(43) <= signed(10,data_width);
      all_coeffs(44) <= signed(10,data_width);
      all_coeffs(45) <= signed(2,data_width);
      all_coeffs(46) <= signed(11,data_width);
      all_coeffs(47) <= signed(5,data_width);
      all_coeffs(48) <= signed(11,data_width);
      all_coeffs(49) <= signed(3,data_width);
      all_coeffs(50) <= signed(13,data_width);
      all_coeffs(51) <= signed(13,data_width);
      all_coeffs(52) <= signed(8,data_width);
      all_coeffs(53) <= signed(8,data_width);
      all_coeffs(54) <= signed(8,data_width);
      all_coeffs(55) <= signed(1,data_width);
      all_coeffs(56) <= signed(6,data_width);
      all_coeffs(57) <= signed(6,data_width);
      all_coeffs(58) <= signed(15,data_width);
      all_coeffs(59) <= signed(12,data_width);
      all_coeffs(60) <= signed(12,data_width);
      all_coeffs(61) <= signed(4,data_width);
      all_coeffs(62) <= signed(9,data_width);
      all_coeffs(63) <= signed(12,data_width);
      all_coeffs(64) <= signed(2,data_width);
      all_coeffs(65) <= signed(13,data_width);
      all_coeffs(66) <= signed(4,data_width);
      all_coeffs(67) <= signed(14,data_width);
      all_coeffs(68) <= signed(10,data_width);
      all_coeffs(69) <= signed(0,data_width);
      all_coeffs(70) <= signed(4,data_width);
      all_coeffs(71) <= signed(4,data_width);
      all_coeffs(72) <= signed(13,data_width);
      all_coeffs(73) <= signed(8,data_width);
      all_coeffs(74) <= signed(14,data_width);
      all_coeffs(75) <= signed(9,data_width);
      all_coeffs(76) <= signed(1,data_width);
      all_coeffs(77) <= signed(8,data_width);
      all_coeffs(78) <= signed(12,data_width);
      all_coeffs(79) <= signed(2,data_width);
      all_coeffs(80) <= signed(7,data_width);
      all_coeffs(81) <= signed(10,data_width);
      all_coeffs(82) <= signed(8,data_width);
      all_coeffs(83) <= signed(3,data_width);
      all_coeffs(84) <= signed(14,data_width);
      all_coeffs(85) <= signed(2,data_width);
      all_coeffs(86) <= signed(4,data_width);
      all_coeffs(87) <= signed(0,data_width);
      all_coeffs(88) <= signed(15,data_width);
      all_coeffs(89) <= signed(15,data_width);
      all_coeffs(90) <= signed(11,data_width);
      all_coeffs(91) <= signed(6,data_width);
      all_coeffs(92) <= signed(10,data_width);
      all_coeffs(93) <= signed(11,data_width);
      all_coeffs(94) <= signed(14,data_width);
      all_coeffs(95) <= signed(4,data_width);
      all_coeffs(96) <= signed(9,data_width);
      all_coeffs(97) <= signed(10,data_width);
      all_coeffs(98) <= signed(6,data_width);
      all_coeffs(99) <= signed(15,data_width);
      all_coeffs(100) <= signed(10,data_width);
      all_coeffs(101) <= signed(0,data_width);
      all_coeffs(102) <= signed(12,data_width);
      all_coeffs(103) <= signed(2,data_width);
      all_coeffs(104) <= signed(14,data_width);
      all_coeffs(105) <= signed(5,data_width);
      all_coeffs(106) <= signed(12,data_width);
      all_coeffs(107) <= signed(7,data_width);
      all_coeffs(108) <= signed(11,data_width);
      all_coeffs(109) <= signed(7,data_width);
      all_coeffs(110) <= signed(2,data_width);
      all_coeffs(111) <= signed(0,data_width);
      all_coeffs(112) <= signed(4,data_width);
      all_coeffs(113) <= signed(12,data_width);
      all_coeffs(114) <= signed(1,data_width);
      all_coeffs(115) <= signed(15,data_width);
      all_coeffs(116) <= signed(3,data_width);
      all_coeffs(117) <= signed(12,data_width);
      all_coeffs(118) <= signed(0,data_width);
      all_coeffs(119) <= signed(11,data_width);
      all_coeffs(120)<=signed(1, data_width);
      all_coeffs(121)<=signed(3, data_width);
      all_coeffs(122)<=signed(5, data_width);
      all_coeffs(123)<=signed(1, data_width);
      all_coeffs(124)<=signed(6, data_width);
      all_coeffs(125)<=signed(4, data_width);
      all_coeffs(126)<=signed(2, data_width);
      all_coeffs(127)<=signed(10, data_width);
      all_coeffs(128)<=signed(0, data_width);
      all_coeffs(129)<=signed(2, data_width);
      all_coeffs(130)<=signed(0, data_width);
      all_coeffs(131)<=signed(8, data_width);
      
      --more coefficients to be added
      
      data_out <= all_coeffs(to_integer(rd_addr)); 
END behavior;