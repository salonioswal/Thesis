Library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mypackage2.all;

entity mac is
	
	port (Q0 : in signed (data_width-1 downto 0);
		  Q1 : in signed (data_width-1 downto 0);
		  clock: in std_logic;
		  reset: in std_logic;
		  acc: out signed(2*data_width-1 downto 0);
		  mac_en: in std_logic);
	end mac;
	
architecture behavioral_mac of mac is
	signal reg: signed(2*data_width-1 downto 0):=(OTHERS => '0');
	
begin	
process(clock,reset)
begin
if(reset='0') then
	reg<=(OTHERS => '0');
elsif(rising_edge(clock) and mac_en='1') then
	reg<= Q0*Q1 + reg;
end if;
end process;
acc<= reg;

end behavioral_mac;
