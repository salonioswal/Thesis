library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.my_package.all; 
use work.all;

entity test_Be is
	end test_Be;
	
architecture test_b of test_Be is
	signal data_input		: signed(data_width-1 downto 0);
	signal clock			: std_logic;
	signal reset			: std_logic;
	signal column_counter		: unsigned(ptr_width_inv-1 downto 0);
	signal row_counter		: unsigned(ptr_width_inv-1 downto 0);
	signal mac_en			: std_logic;
	signal mac_reset		: std_logic;
	signal addr	:unsigned(ptr_width_inv-1 downto 0);
	constant time_delay : time := 10 ns;

begin
dut: entity work.BE_inverse
	port map(data_input=>data_input,	
		 clock=>clock,
		 reset=>reset,		
		 column_counter=>column_counter,	
		 row_counter=>row_counter,	
		 mac_en=>mac_en,		
		mac_reset=>mac_reset,
		addr=>addr);
	
simulation: process
begin	addr<="00";
	data_input<=x"0000";
	column_counter<=(others=>'0');
	row_counter<=(others=>'0');
	mac_reset<='1';
	reset<='0';
	mac_en<='1';
	wait for time_delay;
	addr<="00";
	data_input<=x"0001";
	mac_reset<='1';
	reset<='1';
	mac_en<='1';
	wait for time_delay;
	addr<="01";
	data_input<=x"0000";
	wait for time_delay;
	addr<="10";
	data_input<=x"0000";
	wait for time_delay;
	row_counter<="01";
mac_reset<='0';

wait for time_delay;
mac_reset<='1';
mac_en<='1';
	addr<="00";
	data_input<=x"0002";	
	wait for time_delay;
	addr<="01";
	data_input<=x"0001";
	wait for time_delay;
addr<="10";
	data_input<=x"0000";
	wait for time_delay;
	row_counter<="10";
mac_reset<='0';

wait for time_delay;
mac_en<='1';
mac_reset<='1';
addr<="00";

	data_input<=x"0003";	
	wait for time_delay;
addr<="01";
data_input<=x"0007";
	wait for time_delay;
addr<="10";
	data_input<=x"0001";
	wait for time_delay;
	mac_en<='0';
	wait for time_delay;
	wait for time_delay;
end process;	

clkgeneration_FC: process
	begin
		clock<= '1';
		wait for time_delay/2;
		clock<= '0';
	        wait for time_delay/2;
	end process clkgeneration_FC;
				
end test_b;


	



		 			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 