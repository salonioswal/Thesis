library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mypackage2.all; 

entity testbench_conv is
	end testbench_conv;

architecture behv_test of testbench_conv is

signal data_input:  signed(data_width-1 downto 0);
signal data_output:  signed(2*data_width-1 downto 0);
signal clock:  std_logic;
signal sys_reset:  std_logic:='0';
signal reset_shifter: std_logic:='0';
signal reset_mac:  std_logic:='0';
signal wr_ptr:  unsigned (1 downto 0):=(others=>'0');
signal wr_en:  std_logic:='0';
signal rd_ptr:  unsigned (1 downto 0):=(others=>'0');
signal mac_en:  std_logic:='0';
		
constant time_delay : time := 10 ns;
begin
dut: entity work.final_conv

port map(data_input=>data_input,
		 data_output=>data_output,
		 clock=>clock,
		 sys_reset=> sys_reset,
		 reset_shifter=>reset_shifter,
		 reset_mac=>reset_mac,
		 wr_ptr=>wr_ptr,
		 wr_en=>wr_en,
		 rd_ptr=>rd_ptr,
		 mac_en=>mac_en);
	
simulation: process
begin
	data_input<=x"0000";
	sys_reset<='1';
	reset_mac<='1';
	reset_shifter<='1';
	wr_en<= '1';
	wait for time_delay;
	data_input<=x"0000";
	wait for time_delay;
	data_input<=x"0001";
	wr_ptr<="01";
	wait for time_delay;
	data_input<=x"0002";
	wr_ptr<="10";
	wait for time_delay;
	data_input<=x"0003";
	wr_ptr<="11";
	wait for time_delay;
	wr_en<= '0';
	mac_en<='1';
	rd_ptr<="00";
	wait for time_delay;
	rd_ptr<="01";
	wait for time_delay;
	rd_ptr<="10";
	wait for time_delay;
	rd_ptr<="11";
	wait for 4*time_delay;	
end process;	

clkgeneration_FC: process
	begin
		clock<= '1';
		wait for time_delay/2;
		clock<= '0';
	        wait for time_delay/2;
	end process clkgeneration_FC;
				
end behv_test;


	



		 