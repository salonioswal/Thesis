library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.my_package.all; 
use work.all;

entity test_ben is
	end test_ben;

architecture test_beh of test_ben is
	signal input_data: signed(data_width-1 downto 0);
	signal output_data:  m_file;
	signal clock: std_logic;
	signal reset: std_logic:='0';
	signal start: std_logic:='0';
	constant time_delay : time := 10 ns;

begin
dut: entity work.comb_strassen 
	port map(input_data=>input_data,
		 output_data=>output_data,
		 clock=>clock,
		 reset=>reset,
		 start=>start);
	
simulation: process
	begin
	reset<='0';
	wait for time_delay;
	input_data<=x"0000";
	reset<='1';
	start<='1';
	wait for time_delay;
	wait for time_delay;
	input_data<=x"0000";
	wait for time_delay;
	input_data<=x"0001";
	wait for time_delay;
	input_data<=x"0001";
	wait for time_delay;
	input_data<=x"0000";
	wait for time_delay;
	input_data<=x"0000";
	wait for time_delay;
	input_data<=x"0001";
	wait for time_delay;
	input_data<=x"0001";
	wait for time_delay;
	input_data<=x"0000";
	wait for 200*time_delay;
end process;
	
clkgeneration_FC: process
	begin
		clock<= '1';
		wait for time_delay/2;
		clock<= '0';
	        wait for time_delay/2;
	end process clkgeneration_FC;
		
end test_beh;		
		
		
		
		
		
		
		